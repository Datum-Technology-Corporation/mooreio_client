// Copyright 2024 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_MAPU_B_TDEFS_SV__
`define __UVMT_MAPU_B_TDEFS_SV__


// pragma uvmx tdefs begin
// Add enums and structs here
// Ex: typedef bit [(`UVMT_MAPU_B_ABC-1):0]  uvmt_mapu_b_abc_b_t; ///< Describe me!
// Ex: /*
//      * Describe me!
//      */
//     typedef enum {
//        UVMT_MAPU_B_EX_ABC
//     } uvmt_mapu_b_ex_enum;
// Ex: /*
//      * Describe me!
//      */
//     typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_mapu_b_ex_struct;
// pragma uvmx tdefs end


`endif // __UVMT_MAPU_B_TDEFS_SV__
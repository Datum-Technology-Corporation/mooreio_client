// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_MPB_ST_MACROS_SVH__
`define __UVMT_MPB_ST_MACROS_SVH__


`ifndef UVMT_MPB_ST_DATA_WIDTH
   `define UVMT_MPB_ST_DATA_WIDTH 32
`endif
`ifndef UVMT_MPB_ST_ADDR_WIDTH
   `define UVMT_MPB_ST_ADDR_WIDTH 32
`endif

// pragma uvmx macros begin
// pragma uvmx macros end


`endif // __UVMT_MPB_ST_MACROS_SVH__
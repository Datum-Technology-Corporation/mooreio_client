// Copyright 2024 Datron Limited Partnership
// SPDX-License-Identifier: MIT
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MAPU_B_CONSTANTS_SV__
`define __UVMA_MAPU_B_CONSTANTS_SV__


const int unsigned  uvma_mapu_b_default_data_width = 32; ///< Default Data Width


// pragma uvmx constants begin
// pragma uvmx constants end


`endif // __UVMA_MAPU_B_CONSTANTS_SV__
// Copyright 2024 Datron Limited Partnership
// SPDX-License-Identifier: MIT
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MAPU_B_MACROS_SVH__
`define __UVMA_MAPU_B_MACROS_SVH__


`define UVMA_MAPU_B_DATA_WIDTH_MIN  32
`define UVMA_MAPU_B_DATA_WIDTH_MAX  64

// pragma uvmx macros begin
// pragma uvmx macros end


`endif // __UVMA_MAPU_B_MACROS_SVH__
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "tb_macros.svh"


package tb_pkg;
  `include "smoke_test.sv"
endpackage

`include "tb.sv"

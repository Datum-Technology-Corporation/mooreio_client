// Copyright 2023 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __MTX_MACROS_SVH__
`define __MTX_MACROS_SVH__




`endif // __MTX_MACROS_SVH__
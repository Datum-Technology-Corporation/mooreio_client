// Copyright 2024 Datron Limited Partnership
// SPDX-License-Identifier: MIT
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MAPU_B_FTDECS_SV__
`define __UVMA_MAPU_B_FTDECS_SV__


typedef class uvma_mapu_b_cfg_c;
typedef class uvma_mapu_b_cntxt_c;
typedef class uvma_mapu_b_dpi_seq_item_c;
typedef class uvma_mapu_b_dpo_seq_item_c;
typedef class uvma_mapu_b_cp_seq_item_c;
typedef class uvma_mapu_b_idle_drv_seq_c;
typedef class uvma_mapu_b_seq_item_c;
typedef class uvma_mapu_b_mon_seq_c;
typedef class uvma_mapu_b_in_drv_seq_c;
typedef class uvma_mapu_b_out_drv_seq_c;


// pragma uvmx ftdecs begin
// pragma uvmx ftdecs end


`endif // __UVMA_MAPU_B_FTDECS_SV__
import uvm_pkg::*;
`include "uvm_macros.svh"


package def_ss_tb_pkg;
  import uvm_pkg::*;
  `include "def_ss_tb_macros.svh"
  `include "def_ss_smoke_test.sv"
endpackage

`include "def_ss_tb.sv"

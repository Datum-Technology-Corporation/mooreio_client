// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_MPB_ST_FTDECS_SV__
`define __UVMT_MPB_ST_FTDECS_SV__


// pragma uvmx ftdecs begin
// pragma uvmx ftdecs end


`endif // __UVMT_MPB_ST_FTDECS_SV__
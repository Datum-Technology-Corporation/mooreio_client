// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_MAPU_B_BASE_TEST_WORKAROUNDS_SV__
`define __UVMT_MAPU_B_BASE_TEST_WORKAROUNDS_SV__


// pragma uvmx base_test_workarounds begin
// Temporary configuration constraints belong here (this file should be empty by the end of the project).
// pragma uvmx base_test_workarounds end


`endif // __UVMT_MAPU_B_BASE_TEST_WORKAROUNDS_SV__
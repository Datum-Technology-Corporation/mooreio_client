// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MSTREAM_MACROS_SVH__
`define __UVMA_MSTREAM_MACROS_SVH__


`define UVMA_MSTREAM_DATA_WIDTH_MIN  32
`define UVMA_MSTREAM_DATA_WIDTH_MAX  64

// pragma uvmx macros begin
// pragma uvmx macros end


`endif // __UVMA_MSTREAM_MACROS_SVH__
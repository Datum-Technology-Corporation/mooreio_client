// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MAPU_B_IF_CHKR_SV__
`define __UVMA_MAPU_B_IF_CHKR_SV__


/**
 * Module encapsulating assertions targeting Matrix APU Block Agent interface.
 * @ingroup uvma_mapu_b_pkg
 */
module uvma_mapu_b_if_chkr (
   uvma_mapu_b_if  agent_if ///< Target interface
);

   // pragma uvmx interface_checker begin
   // pragma uvmx interface_checker end

endmodule


`endif // __UVMA_MAPU_B_IF_CHKR_SV__
// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MSTREAM_ST_FTDECS_SV__
`define __UVME_MSTREAM_ST_FTDECS_SV__


typedef class uvme_mstream_st_base_seq_c;
typedef class uvme_mstream_st_fix_stim_seq_c;
typedef class uvme_mstream_st_rand_stim_seq_c;

// pragma uvmx ftdecs begin
// pragma uvmx ftdecs end


`endif // __UVME_MSTREAM_ST_FTDECS_SV__
module block_top();

endmodule : block_top
// Copyright 2024 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MAPU_B_CONSTANTS_SV__
`define __UVME_MAPU_B_CONSTANTS_SV__


// pragma uvmx constants begin
// pragma uvmx constants end


`endif // __UVME_MAPU_B_CONSTANTS_SV__
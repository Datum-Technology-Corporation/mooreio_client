// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MSTREAM_FTDECS_SV__
`define __UVMA_MSTREAM_FTDECS_SV__


typedef class uvma_mstream_cfg_c;
typedef class uvma_mstream_cntxt_c;
typedef class uvma_mstream_pkt_seq_item_c;
typedef class uvma_mstream_pkt_mon_trn_c;
typedef class uvma_mstream_host_ig_seq_item_c;
typedef class uvma_mstream_card_ig_seq_item_c;
typedef class uvma_mstream_ig_mon_trn_c;
typedef class uvma_mstream_host_eg_seq_item_c;
typedef class uvma_mstream_card_eg_seq_item_c;
typedef class uvma_mstream_eg_mon_trn_c;
typedef class uvma_mstream_ig_mon_seq_c;
typedef class uvma_mstream_eg_mon_seq_c;
typedef class uvma_mstream_idle_drv_seq_c;
typedef class uvma_mstream_pkt_drv_seq_c;
typedef class uvma_mstream_rx_drv_seq_c;
typedef class uvma_mstream_pkt_base_seq_c;
typedef class uvma_mstream_pkt_rand_stim_seq_c;

// pragma uvmx ftdecs begin
// pragma uvmx ftdecs end


`endif // __UVMA_MSTREAM_FTDECS_SV__
// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MAPU_B_ENV_SV__
`define __UVME_MAPU_B_ENV_SV__


/**
 * Matrix APU Block UVM Environment with TLM prediction.
 * @ingroup uvme_mapu_b_comps
 */
class uvme_mapu_b_env_c extends uvmx_block_env_c #(
   .T_CFG      (uvme_mapu_b_cfg_c      ),
   .T_CNTXT    (uvme_mapu_b_cntxt_c    ),
   .T_SQR      (uvme_mapu_b_sqr_c      ),
   .T_PRD      (uvme_mapu_b_prd_c      ),
   .T_SB       (uvme_mapu_b_sb_c       ),
   .T_COV_MODEL(uvme_mapu_b_cov_model_c)
);

   /// @name Agents
   /// @{
   uvma_mapu_b_agent_c  agent; ///< Block agent
   /// @}

   /// @name Ports
   /// @{
   uvm_analysis_port #(uvma_mapu_b_ig_mon_trn_c)  monitored_ig_ap; ///< Monitored ingress
   uvm_analysis_port #(uvma_mapu_b_eg_mon_trn_c)  monitored_eg_ap; ///< Monitored egress
   uvm_analysis_port #(uvma_mapu_b_eg_mon_trn_c)  predicted_eg_ap; ///< Predicted egress
   /// @}

   // pragma uvmx env_fields begin
   // pragma uvmx env_fields end


   `uvm_component_utils_begin(uvme_mapu_b_env_c)
      // pragma uvmx env_uvm_field_macros begin
      // pragma uvmx env_uvm_field_macros end
   `uvm_component_utils_end


   /**
    * Default constructor.
    */
   function new(string name="uvme_mapu_b_env", uvm_component parent=null);
      super.new(name, parent);
   endfunction

   /**
    * Assigns configuration handles to components using UVM Configuration Database.
    */
   virtual function void assign_cfg();
      uvm_config_db#(uvma_mapu_b_cfg_c)::set(this, "agent", "cfg", cfg.agent_cfg);
      // pragma uvmx env_assign_cfg begin
      // pragma uvmx env_assign_cfg end
   endfunction

   /**
    * Assigns context handles to components using UVM Configuration Database.
    */
   virtual function void assign_cntxt();
      uvm_config_db#(uvma_mapu_b_cntxt_c)::set(this, "agent", "cntxt", cntxt.agent_cntxt);
      // pragma uvmx env_assign_cntxt begin
      // pragma uvmx env_assign_cntxt end
   endfunction

   /**
    * Creates agent components.
    */
   virtual function void create_agents();
      agent = uvma_mapu_b_agent_c::type_id::create("agent", this);
      // pragma uvmx env_create_agents begin
      // pragma uvmx env_create_agents end
   endfunction

   /**
    * Connects agents to predictor.
    */
   virtual function void connect_predictor();
      agent.ig_mon_trn_ap.connect(predictor.ig_fifo.analysis_export);
      // pragma uvmx env_connect_predictor begin
      // pragma uvmx env_connect_predictor end
   endfunction

   /**
    * Connects scoreboards components to agents/predictor.
    */
   virtual function void connect_scoreboard();
      predictor.eg_ap.connect(scoreboard.egress_scoreboard.exp_export);
      agent.eg_mon_trn_ap.connect(scoreboard.egress_scoreboard.act_export);
      // pragma uvmx env_connect_scoreboard begin
      // pragma uvmx env_connect_scoreboard end
   endfunction

   /**
    * Connects environment coverage model to agent/predictor.
    */
   virtual function void connect_coverage_model();
      agent.seq_item_ap.connect(cov_model.agent_op_fifo.analysis_export);
      agent.ig_mon_trn_ap.connect(cov_model.agent_ig_fifo.analysis_export);
      predictor.eg_ap.connect(cov_model.predictor_eg_fifo.analysis_export);
      agent.cp_seq_item_ap.connect(cov_model.agent_cp_stim_fifo.analysis_export);
      agent.cp_mon_trn_ap.connect(cov_model.agent_cp_mon_fifo.analysis_export);
      // pragma uvmx env_connect_coverage_model begin
      // pragma uvmx env_connect_coverage_model end
   endfunction

   /**
    * Connects environment output ports to components.
    */
   virtual function void connect_ports();
      monitored_ig_ap = agent.ig_mon_trn_ap;
      monitored_eg_ap = agent.eg_mon_trn_ap;
      predicted_eg_ap = predictor.eg_ap;
      // pragma uvmx env_connect_ports begin
      // pragma uvmx env_connect_ports end
   endfunction

   /**
    * Assembles sequencer from agent sequencers.
    */
   virtual function void assemble_sequencer();
      sequencer.agent_sequencer = agent.sequencer;
      // pragma uvmx env_start_sequences begin
      // pragma uvmx env_start_sequences end
   endfunction

   // pragma uvmx env_methods begin
   // pragma uvmx env_methods end

endclass


`endif // __UVME_MAPU_B_ENV_SV__
// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_MPB_ST_TDEFS_SV__
`define __UVMT_MPB_ST_TDEFS_SV__


// pragma uvmx tdefs begin
// Add enums and structs here
// Ex: typedef bit [(`UVMT_MPB_ST_ABC-1):0]  uvmt_mpb_st_abc_b_t; ///< Describe me!
// Ex: /*
//      * Describe me!
//      */
//     typedef enum {
//        UVMT_MPB_ST_EX_ABC
//     } uvmt_mpb_st_ex_enum;
// Ex: /*
//      * Describe me!
//      */
//     typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_mpb_st_ex_struct;
// pragma uvmx tdefs end


`endif // __UVMT_MPB_ST_TDEFS_SV__
// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MSTREAM_ST_CONSTANTS_SV__
`define __UVME_MSTREAM_ST_CONSTANTS_SV__


// pragma uvmx constants begin
// pragma uvmx constants end


`endif // __UVME_MSTREAM_ST_CONSTANTS_SV__
// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MAPU_B_FTDECS_SV__
`define __UVME_MAPU_B_FTDECS_SV__


// pragma uvmx ftdecs begin
// pragma uvmx ftdecs end


`endif // __UVME_MAPU_B_FTDECS_SV__
// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MSTREAM_CONSTANTS_SV__
`define __UVMA_MSTREAM_CONSTANTS_SV__


const int unsigned  uvma_mstream_default_data_width = 32; ///< Default Data Width


// pragma uvmx constants begin
// pragma uvmx constants end


`endif // __UVMA_MSTREAM_CONSTANTS_SV__
// Copyright 2024 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MAPU_B_MACROS_SVH__
`define __UVME_MAPU_B_MACROS_SVH__


// pragma uvmx macros begin
// Add preprocessor macros here
// Ex: `ifndef UVME_MAPU_B_ABC
//        `define UVME_MAPU_B_ABC 32
//     `endif
// pragma uvmx macros end


`endif // __UVME_MAPU_B_MACROS_SVH__
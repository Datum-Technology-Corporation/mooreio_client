module ss_top();
    block_top  block_instance();
endmodule : ss_top
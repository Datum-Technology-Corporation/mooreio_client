// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MPB_CONSTANTS_SV__
`define __UVMA_MPB_CONSTANTS_SV__


const int unsigned  uvma_mpb_default_data_width = 32; ///< Default Data Width
const int unsigned  uvma_mpb_default_addr_width = 32; ///< Default Address Width


// pragma uvmx constants begin
// pragma uvmx constants end


`endif // __UVMA_MPB_CONSTANTS_SV__
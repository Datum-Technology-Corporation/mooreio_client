module def_ss_top #(
  parameter DATA_WIDTH=8
) (
  input    clk,
  input  rst_n,
  output [(DATA_WIDTH-1):0] o_data_0,
  output [(DATA_WIDTH-1):0] o_data_1
);
endmodule

// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MPB_ST_MACROS_SVH__
`define __UVME_MPB_St_MACROS_SVH__


// pragma uvmx macros begin
// Add preprocessor macros here
// Ex: `ifndef UVME_MPB_ST_ABC
//        `define UVME_MPB_ST_ABC 32
//     `endif
// pragma uvmx macros end


`endif // __UVME_MPB_ST_MACROS_SVH__
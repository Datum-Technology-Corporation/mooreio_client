// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_MAPU_B_MACROS_SVH__
`define __UVMT_MAPU_B_MACROS_SVH__


`ifndef UVMT_MAPU_B_DATA_WIDTH
   `define UVMT_MAPU_B_DATA_WIDTH 32
`endif

// pragma uvmx macros begin
// pragma uvmx macros end


`endif // __UVMT_MAPU_B_MACROS_SVH__
// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MAPU_B_FTDECS_SV__
`define __UVME_MAPU_B_FTDECS_SV__


typedef class uvme_mapu_b_base_seq_c;
typedef class uvme_mapu_b_fix_stim_seq_c;
typedef class uvme_mapu_b_fix_ill_stim_seq_c;
typedef class uvme_mapu_b_rand_stim_seq_c;
typedef class uvme_mapu_b_rand_ill_stim_seq_c;

// pragma uvmx ftdecs begin
// pragma uvmx ftdecs end


`endif // __UVME_MAPU_B_FTDECS_SV__
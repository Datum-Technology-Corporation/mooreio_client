// Copyright 2025 Datron Limited Partnership
// SPDX-License-Identifier: MIT
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MPB_FTDECS_SV__
`define __UVMA_MPB_FTDECS_SV__


typedef class uvma_mpb_cfg_c;
typedef class uvma_mpb_cntxt_c;
typedef class uvma_mpb_access_seq_item_c;
typedef class uvma_mpb_access_mon_trn_c;
typedef class uvma_mpb_main_p_seq_item_c;
typedef class uvma_mpb_sec_p_seq_item_c;
typedef class uvma_mpb_p_mon_trn_c;
typedef class uvma_mpb_access_mon_seq_c;
typedef class uvma_mpb_idle_drv_seq_c;
typedef class uvma_mpb_access_drv_seq_c;
typedef class uvma_mpb_rsp_drv_seq_c;
typedef class uvma_mpb_rsp_base_seq_c;
typedef class uvma_mpb_rsp_mem_seq_c;

// pragma uvmx ftdecs begin
// pragma uvmx ftdecs end


`endif // __UVMA_MPB_FTDECS_SV__